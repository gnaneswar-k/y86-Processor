module ALU_64_2_tb;

parameter WIDTH = 64; //-9223372036854775808 to +9223372036854775807

reg [1:0] S;
reg signed [WIDTH - 1:0] A, B;
wire signed [WIDTH - 1:0] Y;
wire OF;

ALU_64_2 ALU(.Y(Y),.A(A),.B(B),.S(S),.OF(OF));

initial begin
	$dumpfile("ALU_64_2_tb.vcd");
	$dumpvars(0,ALU_64_2_tb);
	$display("S = 00 --> ADD\nS = 01 --> SUB\nS = 10 --> AND\nS = 11 --> XOR");
	S = 2'd0;
	A = 64'sd0;
	B = 64'sd0;
end

initial begin
	$monitor("time =%0t \t S =%b, A =%0d, B =%0d, Y =%0d, OF =%b",$time,S,A,B,Y,OF);
	S = 2'd0;
	A = 64'sd0;//0
	B = 64'sd0;//0
	
	#10;
	S = 2'd1;
	
	#10;
	S = 2'd2;
	
	#10;
	S = 2'd3;
	
	#10;
	S = 2'd0;
	A = 64'sd1;//1
	B = -64'sd1;//-1
	
	#10;
	S = 2'd1;
	
	#10;
	S = 2'd2;
	
	#10;
	S = 2'd3;
	
	#10;
	S = 2'd0;
	A = 64'sd9223372036854775807;//9223372036854775807
	B = 64'sd9223372036854775807;//9223372036854775807
	
	#10;
	S = 2'd1;
	
	#10;
	S = 2'd2;
	
	#10;
	S = 2'd3;
	
	#10;
	S = 2'd0;
	A = 64'sd9223372036854775807;//9223372036854775807
	B = -64'sd9223372036854775808;//-9223372036854775808
	
	#10;
	S = 2'd1;
	
	#10;
	S = 2'd2;
	
	#10;
	S = 2'd3;
	
	#10;
	S = 2'd0;
	A = 64'sd0;//0;
	B = -64'sd9223372036854775808;//-9223372036854775808
	
	#10;
	S = 2'd1;
	
	#10;
	S = 2'd2;
	
	#10;
	S = 2'd3;
	
	#10;
	S = 2'd0;
	A = -64'sd9223372036854775808;//-9223372036854775808
	B = 64'sd0;//0
	
	#10;
	S = 2'd1;
	
	#10;
	S = 2'd2;
	
	#10;
	S = 2'd3;
	
	#10;
	S = 2'd0;
	A = -64'sd9223372036854775808;//-9223372036854775808
	B = -64'sd9223372036854775808;//-9223372036854775808
	
	#10;
	S = 2'd1;
	
	#10;
	S = 2'd2;
	
	#10;
	S = 2'd3;
	
	#10;
	S = 2'd0;
	A = 64'sd0;//0
	B = 64'sd0;//0
end

endmodule